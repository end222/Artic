-- Author: Pablo Orduna Lagarma
-- Artic Risc V


library ieee;
use ieee.std_logic_1164.all;

entity decode_exec is
	Port (
		in_clk : in std_logic;
		in_reset : in std_logic;
		in_load : in std_logic;

		decode_rs_value : in std_logic_vector(31 downto 0);
		decode_rt_value : in std_logic_vector(31 downto 0);
		decode_rs_id : in std_logic_vector(4 downto 0);
		decode_rt_id : in std_logic_vector(4 downto 0);
		decode_rd_id : in std_logic_vector(4 downto 0);
		decode_inm : in std_logic_vector(31 downto 0);
		decode_rst_inuse : in std_logic; -- Use of RD for risk detection
		decode_fp_add : in std_logic;
		decode_alu_opctrl : in std_logic_vector(1 downto 0);
		decode_memwrite : in std_logic;
		decode_memread : in std_logic;
		-- Determines whether to use ALU output or MEM output to write to the RD reg
		decode_memtoreg : in std_logic;
		-- Determines whether to use inm or RT value 
		decode_alu_src : in std_logic;

		exec_rs_value : out std_logic_vector(31 downto 0);
		exec_rt_value : out std_logic_vector(31 downto 0);
		exec_rs_id : out std_logic_vector(4 downto 0);
		exec_rt_id : out std_logic_vector(4 downto 0);
		exec_rd_id : out std_logic_vector(4 downto 0);
		exec_inm : out std_logic_vector(31 downto 0);
		exec_rst_inuse : out std_logic;
		exec_fp_add : out std_logic;
		exec_alu_opctrl : out std_logic_vector(1 downto 0);
		exec_memwrite : out std_logic;
		exec_memread : out std_logic;
		exec_memtoreg : out std_logic;
		exec_alu_src : out std_logic
	);
end decode_exec;


architecture RTL of decode_exec is
begin
	process(in_clk)
	begin
		if(rising_edge(in_clk)) then
			if (in_reset = '1') then
				exec_rs_value <= "00000000000000000000000000000000";
				exec_rt_value <= "00000000000000000000000000000000";
				exec_rs_id <= "00000";
				exec_rt_id <= "00000";
				exec_rd_id <= "00000";
				exec_inm <= "00000000000000000000000000000000";
				exec_rst_inuse <= '0';
				exec_fp_add <= '0';
				exec_alu_opctrl <= "00";
				exec_memwrite <= '0';
				exec_memread <= '0';
				exec_memtoreg <= '0';
				exec_alu_src <= '0';

			else
				if (in_load = '1') then
					exec_rs_value <= decode_rs_value;
					exec_rt_value <= decode_rt_value;
					exec_rs_id <= decode_rs_id;
					exec_rt_id <= decode_rt_id;
					exec_rd_id <= decode_rd_id;
					exec_inm <= decode_inm;
					exec_rst_inuse <= decode_rst_inuse;
					exec_fp_add <= decode_fp_add;
					exec_alu_opctrl <= decode_alu_opctrl;
					exec_memwrite <= decode_memwrite;
					exec_memread <= decode_memread;
					exec_memtoreg <= decode_memtoreg;
					exec_alu_src <= decode_alu_src;
				end if;
			end if;
		end if;
	end process;
end RTL;
